* SPICE3 file created from BGR.ext - technology: sky130A

.option scale=0.005u

X0 F VBGP VSSA sky130_fd_pr__res_xhigh_po w=70 l=9550
X3 E J VSSA sky130_fd_pr__res_xhigh_po w=70 l=1044
X7 K VDDA VSSA sky130_fd_pr__res_xhigh_po w=70 l=6998

X1 sky130_fd_pr__pnp_05v5_W3p40L3p40_0/c_153_607# VSSA E VSSA sky130_fd_pr__pnp_05v0 area=0
X2 sky130_fd_pr__pnp_05v5_W3p40L3p40_1/c_153_607# VSSA E VSSA sky130_fd_pr__pnp_05v0 area=0
X4 sky130_fd_pr__pnp_05v5_W3p40L3p40_3/c_153_607# VSSA E VSSA sky130_fd_pr__pnp_05v0 area=0
X5 sky130_fd_pr__pnp_05v5_W3p40L3p40_2/c_153_607# VSSA E VSSA sky130_fd_pr__pnp_05v0 area=0
X6 sky130_fd_pr__pnp_05v5_W3p40L3p40_4/c_153_607# VSSA I VSSA sky130_fd_pr__pnp_05v0 area=8.4466e+08
X8 sky130_fd_pr__pnp_05v5_W3p40L3p40_5/c_153_607# VSSA F VSSA sky130_fd_pr__pnp_05v0 area=7
X9 sky130_fd_pr__pnp_05v5_W3p40L3p40_6/c_153_607# VSSA E VSSA sky130_fd_pr__pnp_05v0 area=0
X10 sky130_fd_pr__pnp_05v5_W3p40L3p40_7/c_153_607# VSSA E VSSA sky130_fd_pr__pnp_05v0 area=0
X11 sky130_fd_pr__pnp_05v5_W3p40L3p40_8/c_153_607# VSSA E VSSA sky130_fd_pr__pnp_05v0 area=0
X13 sky130_fd_pr__pnp_05v5_W3p40L3p40_9/c_153_607# VSSA E VSSA  sky130_fd_pr__pnp_05v0 area=0

X12 B En I VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=3137 ps=0 w=4000 l=1000
X14 D A C VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=-1 pd=-1 as=113 ps=0 w=4000 l=1000
X15 A A B VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=4705 pd=0 as=0 ps=0 w=4000 l=1000
X16 J En D VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=3.58118e+06 pd=0 as=-0 ps=-0 w=4000 l=1000
X17 H En VBGP VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=-1 ps=32666 w=4000 l=1000
X18 C G VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=97 ps=0 w=4000 l=1000
X19 G En K VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=86544 pd=0 as=-1 ps=-1 w=4000 l=1000
X20 G A VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=4000 l=200
X21 A C VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=4000 l=1000
X22 C C VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=4000 l=1000
X23 H C VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=4000 l=1000

C0 VBGP En 0.22fF
C1 VBGP C 0.55fF
C2 I A 0.12fF
C3 VDDA A 0.10fF
C4 En A 0.53fF
C5 A G 0.12fF
C6 C A 0.67fF
C7 I J 0.28fF
C8 VDDA C 0.09fF
C9 G K 0.25fF
C10 En G 0.65fF
C11 En C 0.61fF
C12 VDDA H 0.04fF
C13 VBGP A 0.28fF
C14 VBGP K 0.27fF
C15 VDDA VSSA 82.23fF
C16 E VSSA 10.56fF
