* General Purpose Bandgap Reference circuit avsdbgp_3v3- Technology: sky130

.options savecurrents
.lib "/home/anmol/Desktop/vsdflow/work/tools/openlane_working_dir/pdks/skywater-pdk/libraries/sky130_fd_pr/latest/models/sky130.lib.spice" tt
.include "/home/anmol/Desktop/vsdflow/work/tools/openlane_working_dir/pdks/skywater-pdk/libraries/sky130_fd_pr/latest/models/corners/tt/nonfet.spice"
.include "/home/anmol/Desktop/vsdflow/work/tools/openlane_working_dir/pdks/skywater-pdk/libraries/sky130_fd_pr/latest/models/sky130_fd_pr__model__pnp.model.spice"


*BGR circuit

XM1 A C VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 l=5 w=20
XM2 C C VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 l=5 w=20
XM3 VBGP C VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 l=5 w=20
XM4 A A B GND sky130_fd_pr__nfet_g5v0d10v5 l=5 w=20
XM5 C A D GND sky130_fd_pr__nfet_g5v0d10v5 l=5 w=20

X6 GND GND B GND sky130_fd_pr__pnp_05v5_W3p40L3p40 M=1
X7 GND GND E GND sky130_fd_pr__pnp_05v5_W3p40L3p40 M=8
X8 GND GND F GND sky130_fd_pr__pnp_05v5_W3p40L3p40 M=1

*Start-up circuit

XM9 C G GND GND sky130_fd_pr__nfet_g5v0d10v5 l=0.5 w=2
XM10 G A GND GND sky130_fd_pr__nfet_g5v0d10v5 l=0.5 w=10
R1 D E 30K
R2 F VBGP 272K
R3 GND VBGP 100MEG
R4 VPWR G 25K

VDDA VPWR GND DC 3.3V

.dc temp -40 140 0.1

.control
run
plot deriv(v(VBGP))/1.20

.endc

.end

