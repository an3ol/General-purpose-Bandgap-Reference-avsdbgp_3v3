* General Purpose Bandgap Reference circuit avsdbgp_3v3- Technology: sky130

.options savecurrents
.lib "../libs/models/sky130.lib.spice" tt
.include "../libs/models/sky130_fd_pr__model__pnp.model.spice"

*BGR circuit

XM1 A C VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 l=5 w=20
XM2 C C VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 l=5 w=20
XM3 H C VPWR VPWR sky130_fd_pr__pfet_g5v0d10v5 l=5 w=20
XM4 A A B GND sky130_fd_pr__nfet_g5v0d10v5 l=5 w=20
XM5 C A D GND sky130_fd_pr__nfet_g5v0d10v5 l=5 w=20

X6 GND GND I GND sky130_fd_pr__pnp_05v5_W3p40L3p40 M=1
X7 GND GND E GND sky130_fd_pr__pnp_05v5_W3p40L3p40 M=8
X8 GND GND F GND sky130_fd_pr__pnp_05v5_W3p40L3p40 M=1

*Start-up circuit

XM9 C G GND GND sky130_fd_pr__nfet_g5v0d10v5 l=0.5 w=2
XM10 G A GND GND sky130_fd_pr__nfet_g5v0d10v5 l=0.5 w=10

*Enable circuit

XM11 B En Vx GND sky130_fd_pr__nfet_g5v0d10v5 l=0.5 w=4
XM12 D En Vy GND sky130_fd_pr__nfet_g5v0d10v5 l=0.5 w=4
XM13 H En Vz GND sky130_fd_pr__nfet_g5v0d10v5 l=0.5 w=4
XM14 K En G GND sky130_fd_pr__nfet_g5v0d10v5 l=0.5 w=4

R1 J E 30K
R2 F VBGP 272.5K
R3 GND VBGP 100MEG
R4 VPWR Vw 200K

Vsrc Vx I DC 0V
Vsrc1 Vy J DC 0V
Vsrc2 Vz VBGP DC 0V
Vsrc3 Vw K DC 0V

VDDA VPWR GND DC 3.3V
VD En GND DC 3.3V

.dc temp -40 140 0.1

.control
run
plot v(vbgp) v(f) v(vbgp,f)
plot v(VBGP)
.endc

.end
