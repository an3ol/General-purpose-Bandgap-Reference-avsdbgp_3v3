* General Purpose Bandgap Reference circuit avsdbgp_3v3- Technology: sky130
.lib "../../libs/models/sky130.lib.spice" tt
.include "../../libs/models/sky130_fd_pr__model__pnp.model.spice"


.option scale=0.005u

X0 F VBGP VSSA sky130_fd_pr__res_xhigh_po w=70 l=9250
X3 E J VSSA sky130_fd_pr__res_xhigh_po w=70 l=1044
X7 K VDDA VSSA sky130_fd_pr__res_xhigh_po w=70 l=6998

X1 sky130_fd_pr__pnp_05v5_W3p40L3p40_0/c_153_607# VSSA E sky130_fd_pr__pnp_05v5_W3p40L3p40_0/c_153_607# sky130_fd_pr__pnp_05v5_W3p40L3p40 m=1
X2 sky130_fd_pr__pnp_05v5_W3p40L3p40_1/c_153_607# VSSA E sky130_fd_pr__pnp_05v5_W3p40L3p40_1/c_153_607# sky130_fd_pr__pnp_05v5_W3p40L3p40 m=1
X4 sky130_fd_pr__pnp_05v5_W3p40L3p40_3/c_153_607# VSSA E sky130_fd_pr__pnp_05v5_W3p40L3p40_3/c_153_607# sky130_fd_pr__pnp_05v5_W3p40L3p40 m=1
X5 sky130_fd_pr__pnp_05v5_W3p40L3p40_2/c_153_607# VSSA E sky130_fd_pr__pnp_05v5_W3p40L3p40_2/c_153_607# sky130_fd_pr__pnp_05v5_W3p40L3p40 m=1
X6 sky130_fd_pr__pnp_05v5_W3p40L3p40_4/c_153_607# VSSA I sky130_fd_pr__pnp_05v5_W3p40L3p40_4/c_153_607# sky130_fd_pr__pnp_05v5_W3p40L3p40 m=1
X8 sky130_fd_pr__pnp_05v5_W3p40L3p40_5/c_153_607# VSSA F sky130_fd_pr__pnp_05v5_W3p40L3p40_5/c_153_607# sky130_fd_pr__pnp_05v5_W3p40L3p40 m=1
X9 sky130_fd_pr__pnp_05v5_W3p40L3p40_6/c_153_607# VSSA E sky130_fd_pr__pnp_05v5_W3p40L3p40_6/c_153_607# sky130_fd_pr__pnp_05v5_W3p40L3p40 m=1
X10 sky130_fd_pr__pnp_05v5_W3p40L3p40_7/c_153_607# VSSA E sky130_fd_pr__pnp_05v5_W3p40L3p40_7/c_153_607# sky130_fd_pr__pnp_05v5_W3p40L3p40 m=1
X11 sky130_fd_pr__pnp_05v5_W3p40L3p40_8/c_153_607# VSSA E sky130_fd_pr__pnp_05v5_W3p40L3p40_8/c_153_607# sky130_fd_pr__pnp_05v5_W3p40L3p40 m=1
X13 sky130_fd_pr__pnp_05v5_W3p40L3p40_9/c_153_607# VSSA E sky130_fd_pr__pnp_05v5_W3p40L3p40_9/c_153_607# sky130_fd_pr__pnp_05v5_W3p40L3p40 m=1

XM12 B En I VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=3137 ps=0 w=4000 l=1000
XM14 D A C VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=-1 pd=-1 as=113 ps=0 w=4000 l=1000
XM15 A A B VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=4705 pd=0 as=0 ps=0 w=4000 l=1000
XM16 J En D VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=3.58118e+06 pd=0 as=-0 ps=-0 w=4000 l=1000
XM17 H En VBGP VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=-1 ps=32666 w=4000 l=1000
XM18 C G VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=97 ps=0 w=4000 l=1000
XM19 G En K VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=86544 pd=0 as=-1 ps=-1 w=4000 l=1000
XM20 G A VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=4000 l=200
XM21 A C VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=4000 l=1000
XM22 C C VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=4000 l=1000
XM23 H C VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=4000 l=1000


R3 GND VBGP 100MEG

VSS VSSA GND DC 0V
VDD VDDA GND DC 3.3V
VD En GND DC 3.3V

.dc VDD 2 4 0.1

.control
run
plot v(VBGP)
.endc

.end
