magic
tech sky130A
magscale 1 2
timestamp 1615721042
<< nwell >>
rect 11000 2800 17600 3400
<< pwell >>
rect 6612 -10016 18502 -9002
<< mvndiffc >>
rect 7130 -3990 7170 -3930
rect 13240 -4060 13360 -3940
rect 17840 -4060 17960 -3940
rect 6830 -7870 6870 -7810
rect 10640 -7860 10760 -7740
<< mvpdiffc >>
rect 11440 2240 11560 2360
rect 13640 2240 13754 2352
rect 15840 2240 15954 2352
rect 12640 -1560 12760 -1440
rect 14840 -1560 14960 -1440
rect 17040 -1560 17160 -1440
<< poly >>
rect 11600 -2000 12600 -1700
rect 13800 -2000 14800 -1700
rect 16000 -2000 17000 -1700
rect 11600 -2040 17000 -2000
rect 11600 -2160 11640 -2040
rect 11760 -2160 13640 -2040
rect 13760 -2160 15320 -2040
rect 15440 -2160 17000 -2040
rect 11600 -2200 17000 -2160
rect 7598 -3208 17802 -2800
rect 7600 -3802 8602 -3208
rect 9198 -3640 10198 -3602
rect 9198 -3780 9220 -3640
rect 9380 -3780 10198 -3640
rect 9198 -3804 10198 -3780
rect 10800 -3804 11802 -3208
rect 15198 -3802 16200 -3208
rect 16798 -3802 17800 -3208
rect 6900 -8200 7100 -8002
rect 12200 -8200 13202 -8000
rect 13800 -8200 14800 -8000
rect 6898 -8240 14800 -8200
rect 6898 -8360 13240 -8240
rect 13360 -8360 14800 -8240
rect 6898 -8400 14800 -8360
<< polycont >>
rect 11640 -2160 11760 -2040
rect 13640 -2160 13760 -2040
rect 15320 -2160 15440 -2040
rect 9220 -3780 9380 -3640
rect 13240 -8360 13360 -8240
<< locali >>
rect -1002 2400 -696 2402
rect -1002 2070 -570 2400
rect -1002 686 -894 2070
rect -700 686 -570 2070
rect -1002 396 -570 686
rect 7316 1990 7756 2394
rect 11422 2360 11574 2380
rect 11422 2240 11440 2360
rect 11560 2240 11574 2360
rect 11422 2222 11574 2240
rect 13620 2352 13772 2372
rect 13620 2240 13640 2352
rect 13754 2240 13772 2352
rect 13620 2220 13772 2240
rect 15820 2352 15972 2372
rect 15820 2240 15840 2352
rect 15954 2240 15972 2352
rect 15820 2220 15972 2240
rect 7316 596 7396 1990
rect 7614 596 7756 1990
rect 7316 392 7756 596
rect -1996 -1072 -1498 -406
rect -1996 -2384 -1866 -1072
rect -1612 -2384 -1498 -1072
rect -1996 -3000 -1498 -2384
rect 6702 -884 7222 -390
rect 6702 -2722 6810 -884
rect 7122 -2722 7222 -884
rect 12620 -1440 12780 -1420
rect 12620 -1560 12640 -1440
rect 12760 -1560 12780 -1440
rect 12620 -1580 12780 -1560
rect 14820 -1440 14980 -1420
rect 14820 -1560 14840 -1440
rect 14960 -1560 14980 -1440
rect 14820 -1580 14980 -1560
rect 17020 -1440 17180 -1420
rect 17020 -1560 17040 -1440
rect 17160 -1560 17180 -1440
rect 17020 -1580 17180 -1560
rect 11618 -2040 11780 -2020
rect 11618 -2160 11640 -2040
rect 11760 -2160 11780 -2040
rect 11618 -2182 11780 -2160
rect 13620 -2040 13780 -2020
rect 13620 -2160 13640 -2040
rect 13760 -2160 13780 -2040
rect 13620 -2180 13780 -2160
rect 15300 -2040 15460 -2020
rect 15300 -2160 15320 -2040
rect 15440 -2160 15460 -2040
rect 15300 -2180 15460 -2160
rect 6702 -3008 7222 -2722
rect 9200 -3640 9400 -3620
rect 9200 -3780 9220 -3640
rect 9380 -3780 9400 -3640
rect 9200 -3800 9400 -3780
rect 7110 -3930 7190 -3910
rect 7110 -3990 7130 -3930
rect 7170 -3990 7190 -3930
rect 7110 -4010 7190 -3990
rect 13220 -3940 13380 -3920
rect 13220 -4060 13240 -3940
rect 13360 -4060 13380 -3940
rect 13220 -4080 13380 -4060
rect 17820 -3940 17980 -3920
rect 17820 -4060 17840 -3940
rect 17960 -4060 17980 -3940
rect 17820 -4080 17980 -4060
rect 5396 -4802 6604 -4796
rect 5394 -4936 6604 -4802
rect 5394 -5124 5828 -4936
rect 6166 -5124 6604 -4936
rect 5394 -5226 6604 -5124
rect 5396 -5230 6604 -5226
rect -1248 -6912 -802 -6798
rect -462 -6906 -16 -6792
rect 344 -6906 790 -6792
rect 1142 -6900 1588 -6786
rect -1502 -7460 -1362 -7026
rect -696 -7472 -556 -7038
rect 116 -7460 256 -7026
rect 910 -7456 1050 -7022
rect 1700 -7466 1840 -7032
rect 5404 -7276 6598 -7160
rect 5404 -7514 5624 -7276
rect 6388 -7514 6598 -7276
rect -1260 -7698 -814 -7584
rect -458 -7708 -12 -7594
rect 340 -7698 786 -7584
rect 1146 -7692 1592 -7578
rect 5404 -7600 6598 -7514
rect 10620 -7740 10780 -7720
rect 6806 -7810 6890 -7790
rect 6806 -7870 6830 -7810
rect 6870 -7870 6890 -7810
rect 6806 -7890 6890 -7870
rect 10620 -7860 10640 -7740
rect 10760 -7860 10780 -7740
rect -1508 -8156 -1374 -7988
rect 4980 -8080 5550 -7970
rect -1578 -8230 -1314 -8156
rect -1578 -8306 -1498 -8230
rect -1400 -8306 -1314 -8230
rect -1578 -8356 -1314 -8306
rect 4980 -8302 5130 -8080
rect 5398 -8302 5550 -8080
rect 4980 -8414 5550 -8302
rect 5194 -8640 5360 -8414
rect 10620 -8640 10780 -7860
rect 13220 -8240 13380 -8220
rect 13220 -8360 13240 -8240
rect 13360 -8360 13380 -8240
rect 13220 -8380 13380 -8360
rect 5194 -8800 10780 -8640
rect 5194 -8806 5360 -8800
<< viali >>
rect -894 686 -700 2070
rect 11440 2240 11560 2360
rect 13640 2240 13754 2352
rect 15840 2240 15954 2352
rect 7396 596 7614 1990
rect -1866 -2384 -1612 -1072
rect 6810 -2722 7122 -884
rect 12640 -1560 12760 -1440
rect 14840 -1560 14960 -1440
rect 17040 -1560 17160 -1440
rect 11640 -2160 11760 -2040
rect 13640 -2160 13760 -2040
rect 15320 -2160 15440 -2040
rect 9220 -3780 9380 -3640
rect 7130 -3990 7170 -3930
rect 13240 -4060 13360 -3940
rect 17840 -4060 17960 -3940
rect 5828 -5124 6166 -4936
rect 5624 -7514 6388 -7276
rect 6830 -7870 6870 -7810
rect -1498 -8306 -1400 -8230
rect 5130 -8302 5398 -8080
rect 13240 -8360 13360 -8240
<< metal1 >>
rect -1002 2400 -696 2402
rect -1002 2070 -570 2400
rect 7322 2394 7330 2402
rect -1002 686 -894 2070
rect -700 686 -570 2070
rect -1002 396 -570 686
rect 7308 400 7330 2394
rect 7742 400 7748 2402
rect 11416 2360 11576 2800
rect 11416 2240 11440 2360
rect 11560 2240 11576 2360
rect 11416 2216 11576 2240
rect 13616 2352 13776 2800
rect 13616 2240 13640 2352
rect 13754 2240 13776 2352
rect 13616 2214 13776 2240
rect 15816 2352 15976 2800
rect 15816 2240 15840 2352
rect 15954 2240 15976 2352
rect 15816 2214 15976 2240
rect -1998 -1072 -1518 -396
rect -1998 -2384 -1866 -1072
rect -1612 -2384 -1518 -1072
rect -1998 -3006 -1518 -2384
rect 6702 -884 7222 -390
rect 6702 -2722 6810 -884
rect 7122 -1620 7222 -884
rect 12620 -1440 13380 -1420
rect 9502 -1580 9806 -1534
rect 12620 -1560 12640 -1440
rect 12760 -1560 13380 -1440
rect 12620 -1580 13380 -1560
rect 14820 -1440 15460 -1420
rect 14820 -1560 14840 -1440
rect 14960 -1560 15460 -1440
rect 14820 -1580 15460 -1560
rect 17020 -1440 17980 -1420
rect 17020 -1560 17040 -1440
rect 17160 -1560 17980 -1440
rect 17020 -1580 17980 -1560
rect 9502 -1620 9542 -1580
rect 7122 -1780 9542 -1620
rect 7122 -2722 7222 -1780
rect 9502 -1820 9542 -1780
rect 9760 -1820 9806 -1580
rect 9502 -1858 9806 -1820
rect -1820 -3008 -1596 -3006
rect 6702 -3008 7222 -2722
rect 10220 -2040 11780 -2020
rect 10220 -2160 11640 -2040
rect 11760 -2160 11780 -2040
rect 10220 -2180 11780 -2160
rect -1820 -4900 -1720 -3008
rect 7110 -3640 9400 -3618
rect 7110 -3710 9220 -3640
rect 7110 -3930 7190 -3710
rect 8620 -3780 9220 -3710
rect 9380 -3780 9400 -3640
rect 8620 -3802 9400 -3780
rect 8620 -3924 8780 -3802
rect 10220 -3920 10380 -2180
rect 11618 -2182 11780 -2180
rect 7110 -3990 7130 -3930
rect 7170 -3990 7190 -3930
rect 13220 -3940 13380 -1580
rect 13620 -2040 13780 -2020
rect 13620 -2160 13640 -2040
rect 13760 -2160 13780 -2040
rect 13620 -3920 13780 -2160
rect 15300 -2040 15460 -1580
rect 15300 -2160 15320 -2040
rect 15440 -2160 15460 -2040
rect 15300 -2180 15460 -2160
rect 17820 -3940 17980 -1580
rect 7110 -4010 7190 -3990
rect 13220 -4060 13240 -3940
rect 13360 -4060 13380 -3940
rect 17820 -4060 17840 -3940
rect 17960 -4060 17980 -3940
rect 13220 -4080 13380 -4060
rect 17820 -4080 17980 -4060
rect 5382 -4900 6604 -4802
rect -1820 -4902 -1384 -4900
rect -1820 -5000 -1380 -4902
rect -1480 -5240 -1380 -5000
rect -1476 -6906 -1380 -5240
rect 1720 -4936 6604 -4900
rect 1720 -5020 5828 -4936
rect 1720 -6772 1820 -5020
rect 5380 -5124 5828 -5020
rect 6166 -5124 6604 -4936
rect 5380 -5202 6604 -5124
rect 5394 -5226 6604 -5202
rect -582 -6896 1716 -6804
rect -680 -7600 -582 -6898
rect 5404 -7276 6598 -7160
rect 5404 -7514 5624 -7276
rect 6388 -7514 6598 -7276
rect -1380 -7696 -692 -7604
rect -576 -7696 918 -7598
rect 5404 -7600 6598 -7514
rect 1720 -8118 1820 -7722
rect 6498 -7810 6890 -7790
rect 6498 -7870 6830 -7810
rect 6870 -7870 6890 -7810
rect 6498 -7890 6890 -7870
rect 4980 -8080 5550 -7970
rect 1720 -8120 3386 -8118
rect 4980 -8120 5130 -8080
rect -1578 -8230 -1314 -8156
rect -1578 -8306 -1498 -8230
rect -1400 -8306 -1314 -8230
rect 1720 -8278 5130 -8120
rect 3380 -8280 5130 -8278
rect -1578 -8356 -1314 -8306
rect 4980 -8302 5130 -8280
rect 5398 -8302 5550 -8080
rect -1514 -9000 -1400 -8356
rect 4980 -8414 5550 -8302
rect 6498 -8546 6600 -7890
rect 9018 -8546 9178 -7718
rect 13222 -8220 13384 -7874
rect 13220 -8240 13384 -8220
rect 13220 -8360 13240 -8240
rect 13360 -8360 13384 -8240
rect 13220 -8380 13384 -8360
rect 6500 -9000 6600 -8546
rect 9020 -9000 9178 -8546
rect -3800 -10000 20000 -9000
<< via1 >>
rect -894 686 -700 2070
rect 7330 1990 7742 2402
rect 7330 596 7396 1990
rect 7396 596 7614 1990
rect 7614 596 7742 1990
rect 7330 400 7742 596
rect 9542 -1820 9760 -1580
rect 7440 -4060 7560 -3940
rect 16640 -4060 16760 -3940
rect 5624 -7514 6388 -7276
rect 16240 -7858 16362 -7736
<< metal2 >>
rect -1000 3396 -582 3400
rect -1006 3284 -578 3396
rect -1006 2890 -916 3284
rect -680 2890 -578 3284
rect -1006 2794 -578 2890
rect -900 2408 -696 2794
rect -1006 2400 -696 2408
rect 7254 2402 7796 2416
rect -1006 2380 -570 2400
rect -1002 2070 -570 2380
rect -1002 686 -894 2070
rect -700 686 -570 2070
rect -1002 396 -570 686
rect 7254 400 7330 2402
rect 7742 400 7796 2402
rect 7254 386 7796 400
rect 7404 264 7600 386
rect 7404 182 7606 264
rect 7410 40 7606 182
rect 7420 -3940 7580 40
rect 9546 -1534 9762 3190
rect 9502 -1580 9806 -1534
rect 9502 -1820 9542 -1580
rect 9760 -1820 9806 -1580
rect 9502 -1858 9806 -1820
rect 9560 -2418 9740 -1858
rect 10140 -2418 16100 -2416
rect 9560 -2580 16780 -2418
rect 9560 -2582 10610 -2580
rect 10792 -2582 15540 -2580
rect 7420 -4060 7440 -3940
rect 7560 -4060 7580 -3940
rect 7420 -4080 7580 -4060
rect 16620 -3940 16780 -2580
rect 16620 -4060 16640 -3940
rect 16760 -4060 16780 -3940
rect 16620 -4080 16780 -4060
rect 5404 -7276 6598 -7160
rect 5404 -7514 5624 -7276
rect 6388 -7514 6598 -7276
rect 5404 -7600 6598 -7514
rect 5898 -8302 6100 -7600
rect 5900 -8440 6100 -8302
rect 16220 -7736 16380 -7718
rect 16220 -7858 16240 -7736
rect 16362 -7858 16380 -7736
rect 16220 -8440 16380 -7858
rect 5900 -8600 16380 -8440
<< via2 >>
rect -916 2890 -680 3284
<< metal3 >>
rect -3800 3284 20000 3400
rect -3800 2890 -916 3284
rect -680 2890 20000 3284
rect -3800 2800 20000 2890
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_6
timestamp 1615375237
transform 1 0 -1026 0 1 -7246
box 26 26 770 795
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_5
timestamp 1615375237
transform 1 0 -1824 0 1 -7246
box 26 26 770 795
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_1
timestamp 1615375237
transform 1 0 -1026 0 1 -8046
box 26 26 770 795
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_0
timestamp 1615375237
transform 1 0 -1826 0 1 -8046
box 26 26 770 795
use sub2vsscontact  sub2vsscontact_9
timestamp 1615639835
transform 1 0 -1802 0 1 -10002
box 0 0 400 1000
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_7
timestamp 1615375237
transform 1 0 -226 0 1 -7246
box 26 26 770 795
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_2
timestamp 1615375237
transform 1 0 -226 0 1 -8046
box 26 26 770 795
use sub2vsscontact  sub2vsscontact_10
timestamp 1615639835
transform 1 0 -598 0 1 -10004
box 0 0 400 1000
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_9
timestamp 1615375237
transform 1 0 1374 0 1 -7246
box 26 26 770 795
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_8
timestamp 1615375237
transform 1 0 574 0 1 -7248
box 26 26 770 795
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_4
timestamp 1615375237
transform 1 0 1374 0 1 -8046
box 26 26 770 795
use sky130_fd_pr__pnp_05v5_W3p40L3p40  sky130_fd_pr__pnp_05v5_W3p40L3p40_3
timestamp 1615375237
transform 1 0 574 0 1 -8046
box 26 26 770 795
use sub2vsscontact  sub2vsscontact_11
timestamp 1615639835
transform 1 0 600 0 1 -10002
box 0 0 400 1000
use sub2vsscontact  sub2vsscontact_12
timestamp 1615639835
transform 1 0 1798 0 1 -9996
box 0 0 400 1000
use resistor30k  resistor30k_0
timestamp 1615544414
transform 0 1 9804 -1 0 -3598
box 1198 -4400 4002 -3198
use Nmos120  Nmos120_0
timestamp 1615566045
transform 1 0 6800 0 1 -7902
box 0 -100 400 4100
use sub2vsscontact  sub2vsscontact_0
timestamp 1615639835
transform 1 0 6802 0 1 -10002
box 0 0 400 1000
use sub2vsscontact  sub2vsscontact_1
timestamp 1615639835
transform 1 0 8198 0 1 -10004
box 0 0 400 1000
use Nmos520  Nmos520_6
timestamp 1615565174
transform 1 0 5400 0 1 -7902
box 2000 -100 3400 4100
use sub2vsscontact  sub2vsscontact_2
timestamp 1615639835
transform 1 0 9600 0 1 -10002
box 0 0 400 1000
use Nmos520  Nmos520_5
timestamp 1615565174
transform 1 0 6998 0 1 -7904
box 2000 -100 3400 4100
use nmos2metal1  nmos2metal1_8
timestamp 1615594203
transform 1 0 9018 0 1 -7880
box -20 -20 180 160
use sub2vsscontact  sub2vsscontact_3
timestamp 1615639835
transform 1 0 11000 0 1 -10002
box 0 0 400 1000
use Nmos520  Nmos520_0
timestamp 1615565174
transform 1 0 8602 0 1 -7900
box 2000 -100 3400 4100
use sub2vsscontact  sub2vsscontact_4
timestamp 1615639835
transform 1 0 12400 0 1 -10004
box 0 0 400 1000
use Nmos520  Nmos520_1
timestamp 1615565174
transform 1 0 10002 0 1 -7900
box 2000 -100 3400 4100
use sub2vsscontact  sub2vsscontact_5
timestamp 1615639835
transform 1 0 13796 0 1 -10004
box 0 0 400 1000
use Nmos520  Nmos520_2
timestamp 1615565174
transform 1 0 11598 0 1 -7900
box 2000 -100 3400 4100
use nmos2metal1  nmos2metal1_1
timestamp 1615594203
transform 1 0 13222 0 1 -7880
box -20 -20 180 160
use Nmos520  Nmos520_3
timestamp 1615565174
transform 1 0 12998 0 1 -7900
box 2000 -100 3400 4100
use sub2vsscontact  sub2vsscontact_6
timestamp 1615639835
transform 1 0 15200 0 1 -9998
box 0 0 400 1000
use nmos2metal1  nmos2metal1_5
timestamp 1615594203
transform 1 0 16220 0 1 -7878
box -20 -20 180 160
use Nmos520  Nmos520_4
timestamp 1615565174
transform 1 0 14600 0 1 -7900
box 2000 -100 3400 4100
use sub2vsscontact  sub2vsscontact_8
timestamp 1615639835
transform 1 0 18000 0 1 -10000
box 0 0 400 1000
use sub2vsscontact  sub2vsscontact_7
timestamp 1615639835
transform 1 0 16598 0 1 -10000
box 0 0 400 1000
use resistor273k  resistor273k_0
timestamp 1615550117
transform 1 0 -1584 0 1 -3006
box -400 0 8800 2600
use nmos2metal1  nmos2metal1_7
timestamp 1615594203
transform 1 0 7420 0 1 -4080
box -20 -20 180 160
use nmos2metal1  nmos2metal1_3
timestamp 1615594203
transform 1 0 8620 0 1 -4080
box -20 -20 180 160
use nmos2metal1  nmos2metal1_2
timestamp 1615594203
transform 1 0 10220 0 1 -4080
box -20 -20 180 160
use Pmos520  Pmos520_0
timestamp 1615566544
transform 1 0 11400 0 1 -1600
box -400 -400 1800 4400
use nmos2metal1  nmos2metal1_0
timestamp 1615594203
transform 1 0 13620 0 1 -4080
box -20 -20 180 160
use Pmos520  Pmos520_1
timestamp 1615566544
transform 1 0 13600 0 1 -1600
box -400 -400 1800 4400
use Pmos520  Pmos520_2
timestamp 1615566544
transform 1 0 15800 0 1 -1600
box -400 -400 1800 4400
use nmos2metal1  nmos2metal1_4
timestamp 1615594203
transform 1 0 16620 0 1 -4080
box -20 -20 180 160
use resistor200k  resistor200k_0
timestamp 1615546188
transform 1 0 -602 0 1 396
box -400 0 8352 2000
use vddcontact  vddcontact_0
timestamp 1615585694
transform 1 0 11300 0 1 2800
box 0 0 400 600
use vddcontact  vddcontact_1
timestamp 1615585694
transform 1 0 13500 0 1 2800
box 0 0 400 600
use pmossub2vdd  pmossub2vdd_0
timestamp 1615590023
transform 1 0 12300 0 1 2800
box 0 0 400 600
use pmossub2vdd  pmossub2vdd_1
timestamp 1615590023
transform 1 0 14500 0 1 2800
box 0 0 400 600
use vddcontact  vddcontact_2
timestamp 1615585694
transform 1 0 15700 0 1 2800
box 0 0 400 600
use pmossub2vdd  pmossub2vdd_2
timestamp 1615590023
transform 1 0 16700 0 1 2800
box 0 0 400 600
<< labels >>
rlabel metal3 9618 2886 9618 2886 1 VBGP
rlabel poly 15626 -3234 15626 -3234 1 En
rlabel metal3 18646 3076 18646 3076 1 VDDA
rlabel metal1 18950 -9556 18950 -9556 1 VSSA
rlabel poly 12756 -2104 12756 -2104 1 C
rlabel poly 14250 -8280 14250 -8280 1 A
rlabel metal1 17898 -2664 17898 -2664 1 H
rlabel metal2 6000 -8204 6000 -8204 1 J
rlabel metal1 7246 -3668 7246 -3668 1 G
rlabel metal1 3408 -4962 3408 -4962 1 E
rlabel metal1 -1770 -4888 -1770 -4888 1 F
rlabel metal1 2104 -8192 2104 -8192 1 I
rlabel metal1 3012 -9578 3012 -9578 1 VSSA
flabel metal3 18638 3072 18702 3120 0 FreeSans 2400 0 0 0 VDDA
flabel metal1 19126 -9618 19126 -9618 0 FreeSans 2400 0 0 0 VSSA
flabel poly 11152 -3194 11152 -3194 0 FreeSans 1600 0 0 0 En
flabel poly 14342 -2064 14342 -2064 0 FreeSans 1600 0 0 0 C
flabel poly 12592 -8244 12592 -8244 0 FreeSans 1600 0 0 0 A
<< end >>
