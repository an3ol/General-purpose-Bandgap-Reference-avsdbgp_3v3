* SPICE3 file created from BGR.ext - technology: sky130A

.option scale=5000u

X0 F li_6702_n3008# VSSA sky130_fd_pr__res_xhigh_po w=2600 l=8212
X1 E VSSA sky130_fd_pr__pnp_05v5_W3p40L3p40_0/c_153_607# sky130_fd_pr__pnp_05v0 area=112
X2 E VSSA sky130_fd_pr__pnp_05v5_W3p40L3p40_1/c_153_607# sky130_fd_pr__pnp_05v0 area=0
X3 E J VSSA sky130_fd_pr__res_xhigh_po w=1200 l=1928
X4 E VSSA sky130_fd_pr__pnp_05v5_W3p40L3p40_3/c_153_607# sky130_fd_pr__pnp_05v0 area=0
X5 E VSSA sky130_fd_pr__pnp_05v5_W3p40L3p40_2/c_153_607# sky130_fd_pr__pnp_05v0 area=0
X6 I VSSA sky130_fd_pr__pnp_05v5_W3p40L3p40_4/c_153_607# sky130_fd_pr__pnp_05v0 area=0
X7 VDDA li_7316_392# VSSA sky130_fd_pr__res_xhigh_po w=2000 l=7888
X8 F VSSA sky130_fd_pr__pnp_05v5_W3p40L3p40_5/c_153_607# sky130_fd_pr__pnp_05v0 area=0
X9 E VSSA sky130_fd_pr__pnp_05v5_W3p40L3p40_6/c_153_607# sky130_fd_pr__pnp_05v0 area=0
X10 E VSSA sky130_fd_pr__pnp_05v5_W3p40L3p40_7/c_153_607# sky130_fd_pr__pnp_05v0 area=0
X11 E VSSA sky130_fd_pr__pnp_05v5_W3p40L3p40_8/c_153_607# sky130_fd_pr__pnp_05v0 area=0
X12 Nmos520_1/a_2000_0# En I VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=-3.35544e+07 pd=-1 as=740 ps=0 w=4000 l=1000
X13 E VSSA sky130_fd_pr__pnp_05v5_W3p40L3p40_9/c_153_607# sky130_fd_pr__pnp_05v0 area=0
X14 Nmos520_3/a_2000_0# A C VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=16384 pd=0 as=0 ps=8 w=4000 l=1000
X15 A A Nmos520_1/a_2000_0# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=-0 ps=-0 w=4000 l=1000
X16 J En Nmos520_3/a_2000_0# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=4000 l=1000
X17 H En li_6702_n3008# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=2 pd=8 as=2 ps=8 w=4000 l=1000
X18 C G VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=8 w=4000 l=1000
X19 G En li_7316_392# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=-1 pd=32672 as=2 ps=8 w=4000 l=1000
X20 G A VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=-0 pd=0 as=0 ps=0 w=4000 l=200
X21 A C VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=-513 ps=-1 w=4000 l=1000
X22 C C VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=-0 ps=-0 w=4000 l=1000
X23 H C VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=-0 ps=-0 w=4000 l=1000
C0 li_6702_n3008# C 0.55fF
C1 A VDDA 0.10fF
C2 C VDDA 0.09fF
C3 li_6702_n3008# VDDA 0.48fF
C4 A En 0.52fF
C5 I A 0.22fF
C6 En C 0.58fF
C7 En li_6702_n3008# 0.22fF
C8 A C 0.57fF
C9 H VDDA 0.04fF
C10 I J 0.16fF
C11 li_7316_392# li_6702_n3008# 0.27fF
C12 A li_6702_n3008# 0.28fF
C13 G En 0.65fF
C14 G li_7316_392# 0.25fF
C15 G A 0.12fF
C16 E VSSA 7.47fF
C17 F VSSA 0.89fF
C18 VDDA VSSA 83.13fF
C19 I VSSA 1.35fF
