* SPICE3 file created from BGR.ext - technology: sky130A

.option scale=0.005u


.lib "/home/anmol/Desktop/vsdflow/work/tools/openlane_working_dir/pdks/skywater-pdk/libraries/sky130_fd_pr/latest/models/sky130.lib.spice" tt
.include "/home/anmol/Desktop/vsdflow/work/tools/openlane_working_dir/pdks/skywater-pdk/libraries/sky130_fd_pr/latest/models/corners/tt/nonfet.spice"
.include "/home/anmol/Desktop/vsdflow/work/tools/openlane_working_dir/pdks/skywater-pdk/libraries/sky130_fd_pr/latest/models/sky130_fd_pr__model__pnp.model.spice"

X0 F XX VSSA sky130_fd_pr__res_xhigh_po w=2600 l=8212
X3 E J VSSA sky130_fd_pr__res_xhigh_po w=1200 l=1928
X7 VDDA K VSSA sky130_fd_pr__res_xhigh_po w=2000 l=7888

X1 sky130_fd_pr__pnp_05v5_W3p40L3p40_1/c_153_607# VSSA E VSSA sky130_fd_pr__pnp_05v5_W3p40L3p40 M=1
X2 sky130_fd_pr__pnp_05v5_W3p40L3p40_1/c_153_607# VSSA E VSSA sky130_fd_pr__pnp_05v5_W3p40L3p40 M=1
X4 sky130_fd_pr__pnp_05v5_W3p40L3p40_1/c_153_607# VSSA E VSSA sky130_fd_pr__pnp_05v5_W3p40L3p40 M=1
X5 sky130_fd_pr__pnp_05v5_W3p40L3p40_1/c_153_607# VSSA E VSSA sky130_fd_pr__pnp_05v5_W3p40L3p40 M=1
X6 sky130_fd_pr__pnp_05v5_W3p40L3p40_4/c_153_607# VSSA I VSSA sky130_fd_pr__pnp_05v5_W3p40L3p40 M=1
X8 sky130_fd_pr__pnp_05v5_W3p40L3p40_5/c_153_607# VSSA F VSSA sky130_fd_pr__pnp_05v5_W3p40L3p40 M=1
X9 sky130_fd_pr__pnp_05v5_W3p40L3p40_1/c_153_607# VSSA E VSSA sky130_fd_pr__pnp_05v5_W3p40L3p40 M=1
X10 sky130_fd_pr__pnp_05v5_W3p40L3p40_1/c_153_607# VSSA E VSSA sky130_fd_pr__pnp_05v5_W3p40L3p40 M=1
X11 sky130_fd_pr__pnp_05v5_W3p40L3p40_1/c_153_607# VSSA E VSSA sky130_fd_pr__pnp_05v5_W3p40L3p40 M=1
X13 sky130_fd_pr__pnp_05v5_W3p40L3p40_1/c_153_607# VSSA E VSSA sky130_fd_pr__pnp_05v5_W3p40L3p40 M=1

XM12 B En I VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=-0 ps=0 w=4000 l=1000
XM14 D A C VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=1 ps=0 w=4000 l=1000
XM15 A A B VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=-1.22537e+09 pd=22031 as=0 ps=0 w=4000 l=1000
XM16 J En D VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=2 pd=0 as=0 ps=0 w=4000 l=1000
XM17 H En XX VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=8.38861e+06 ps=0 w=4000 l=1000
XM18 C G VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=8.38854e+06 ps=0 w=4000 l=1000
XM19 G En K VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1.0728e+09 pd=0 as=9 ps=0 w=4000 l=1000
XM20 G A VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=4000 l=200
XM21 A C VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=-0 pd=0 as=0 ps=0 w=4000 l=1000
XM22 C C VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=4000 l=1000
XM23 H C VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=4000 l=1000

C0 En XX 0.22fF
C1 G K 0.25fF
C2 C A 0.66fF
C3 En G 0.65fF
C4 En A 0.53fF
C5 En C 0.60fF
C6 I J 0.33fF
C7 XX VDDA 0.48fF
C8 I A 0.12fF
C9 A VDDA 0.10fF
C10 VDDA H 0.04fF
C11 XX A 0.28fF
C12 C VDDA 0.09fF
C13 G A 0.12fF
C14 XX C 0.55fF
C15 XX K 0.27fF
C16 F VSSA 0.68fF
C17 VDDA VSSA 83.13fF
C18 E VSSA 12.04fF



VSS VSSA GND DC 0V
VDD VDDA GND DC 3.3V
VD En GND DC 3.3V

.dc temp -40 140 0.1

.control
run
plot v(VBGP)
.endc

.end
